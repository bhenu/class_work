entity test is
end entity test